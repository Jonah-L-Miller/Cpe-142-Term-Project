module registers(
	input [4:0] read_reg1, read_reg2,
	input [4:0] write_reg,
	input [15:0] write_data, r0,
	input reg_write, reset, write_r0,	
	
	output reg [15:0] read_data1, read_data2
	);
	
	reg [15:0] R [15:0];
	
	always@(*) begin
		if (reset) begin
			R[4'h0] = 16'h 0000;
			R[4'h1] = 16'h 7B18;
			R[4'h2] = 16'h 245B;
			R[4'h3] = 16'h FFFF;
			R[4'h4] = 16'h F0FF;
			R[4'h5] = 16'h 0051;
			R[4'h6] = 16'h 6666;
			R[4'h7] = 16'h 00FF;
			R[4'h8] = 16'h FF88;
			R[4'h9] = 16'h 0000;
			R[4'hA] = 16'h 0000;
			R[4'hB] = 16'h 3099;
			R[4'hC] = 16'h CCCC;
			R[4'hD] = 16'h 0002;
			R[4'hE] = 16'h 0011;
			R[4'hF] = 16'h 0000;
		end
		else if (reg_write)
			R[write_reg] = write_data;
		else if (write_r0)
				R[0] = r0;
		else begin
			read_data1 = R[read_reg1];
			read_data2 = R[read_reg2];
		end
		

	end
endmodule
